// adder4.v
// 4-bit ripple-carry adder built from 1-bit full adders
module adder4(
    input  wire [3:0] a,
    input  wire [3:0] b,
    input  wire       cin,
    output wire [3:0] sum,
    output wire       cout
);
    wire c1, c2, c3;
    full_adder_1bit FA0(.a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(c1));
    full_adder_1bit FA1(.a(a[1]), .b(b[1]), .cin(c1 ), .sum(sum[1]), .cout(c2));
    full_adder_1bit FA2(.a(a[2]), .b(b[2]), .cin(c2 ), .sum(sum[2]), .cout(c3));
    full_adder_1bit FA3(.a(a[3]), .b(b[3]), .cin(c3 ), .sum(sum[3]), .cout(cout));
endmodule